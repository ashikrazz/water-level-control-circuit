CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
1137 88 1917 1028
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1305 184 1418 281
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 163 279 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 R
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44550.8 0
0
13 Logic Switch~
5 160 219 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 Q
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44550.8 1
0
13 Logic Switch~
5 157 150 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 P
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44550.8 2
0
9 Inverter~
13 302 279 0 2 22
0 3 4
0
0 0 112 0
6 74LS04
-21 -19 21 -11
2 A1
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3421 0 0
2
44550.8 3
0
9 Inverter~
13 300 202 0 2 22
0 3 5
0
0 0 112 0
6 74LS04
-21 -19 21 -11
2 A2
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
8157 0 0
2
44550.8 4
0
14 Logic Display~
6 517 283 0 1 2
20 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 R3
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44550.8 5
0
14 Logic Display~
6 518 124 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 R4
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
44550.8 6
0
14 Logic Display~
6 518 207 0 1 2
12 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
7 OutputX
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
44550.8 7
0
8 2-In OR~
219 425 225 0 3 22
0 9 8 6
0
0 0 112 0
6 74LS32
-21 -24 21 -16
2 A5
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4747 0 0
2
44550.8 8
0
5 7415~
219 365 265 0 4 22
0 2 7 4 8
0
0 0 112 0
6 74LS15
-21 -28 21 -20
2 A6
-7 -38 7 -30
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
972 0 0
2
44550.8 9
0
5 7415~
219 367 188 0 4 22
0 2 7 5 9
0
0 0 112 0
6 74LS15
-21 -28 21 -20
2 A7
-7 -38 7 -30
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
3472 0 0
2
44550.8 10
0
13
1 0 2 0 0 8320 0 7 0 0 11 4
518 142
518 143
187 143
187 150
0 1 3 0 0 4096 0 0 4 4 0 2
190 279
287 279
2 3 4 0 0 4224 0 4 10 0 0 4
323 279
332 279
332 274
341 274
0 1 3 0 0 8320 0 0 6 5 0 4
190 279
190 313
517 313
517 301
1 1 3 0 0 0 0 5 1 0 0 4
285 202
202 202
202 279
175 279
2 3 5 0 0 4224 0 5 11 0 0 4
321 202
332 202
332 197
343 197
1 3 6 0 0 4224 0 8 9 0 0 2
518 225
458 225
0 2 7 0 0 8320 0 0 10 10 0 3
219 219
219 265
341 265
0 1 2 0 0 0 0 0 10 11 0 3
234 150
234 256
341 256
1 2 7 0 0 0 0 2 11 0 0 4
172 219
276 219
276 188
343 188
1 1 2 0 0 0 0 3 11 0 0 4
169 150
276 150
276 179
343 179
4 2 8 0 0 4224 0 10 9 0 0 3
386 265
386 234
412 234
4 1 9 0 0 4224 0 11 9 0 0 3
388 188
388 216
412 216
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
6 227 187 251
16 234 176 250
20 Upper Tank Low Sense
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
4 166 193 190
14 174 182 190
21 Upper Tank High Sense
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
7 94 188 118
17 102 177 118
20 Lower Tank Condition
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
518 194 619 218
528 202 608 218
10 Pump Motor
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
467 246 568 270
477 254 557 270
10 Upper Tank
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
471 88 572 112
481 96 561 112
10 Lower Tank
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
